
LIBRARY IEEE;
LIBRARY STD;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;
USE STD.TEXTIO.ALL;


ENTITY M31HDSP200GB180W_4096X8X1CM16 IS 
	PORT (
		CLK	: IN  STD_LOGIC;
		CEN	: IN  STD_LOGIC;
		WEN	: IN  STD_LOGIC;
		A	: IN  STD_LOGIC_VECTOR (11 DOWNTO 0);
		D	: IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		Q	: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
END M31HDSP200GB180W_4096X8X1CM16;

ARCHITECTURE behavioral OF M31HDSP200GB180W_4096X8X1CM16 IS

	TYPE mem_type IS ARRAY (0 TO 4095) OF STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL mem : MEM_TYPE;
	
BEGIN
	
	R_MEM : PROCESS(CLK)	
	BEGIN
		IF CLK = '1' AND CLK'EVENT THEN
			IF CEN = '0' THEN				-- Active Low
				IF WEN = '1' THEN			-- Active Low
					Q <= mem(TO_INTEGER(UNSIGNED(A)));
				END IF;
			END IF;
		END IF;
	END PROCESS;
	
	W_MEM : PROCESS(CLK)	
	BEGIN
		IF CLK = '1' AND CLK'EVENT THEN
			IF CEN = '0' THEN				-- Active Low
				IF WEN = '0' THEN			-- Active Low
					mem(TO_INTEGER(UNSIGNED(A))) <= D;
				END IF;
			END IF;
		END IF;
	END PROCESS;

END behavioral;
	