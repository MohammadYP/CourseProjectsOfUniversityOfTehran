* SPICE netlist written by S-Edit Win32 6.00
* Written on Jan 12, 2025 at 14:45:37

* Waveform probing commands
.probe
.options probefilename="DFlipFlop"
+ probesdbfile="D:\Desktop\Electronic Digital\CA5\part 2\one\DFlipFlop.sdb"
+ probetopmodule="shift_register_4bbit"

* No Ports in cell: PageID_Tanner
* End of module with no ports: PageID_Tanner

.SUBCKT Pad_Bond SIGNAL Subs
C1 SIGNAL Subs 0.25pF
* Page Size:  5x7
* S-Edit  Output Pad
* Designed by: D.Gunawan, J.Luo, K.Schaefer  Jan 12, 2025  14:21:54
* Schematic generated by S-Edit
* from file D:\Desktop\Electronic Digital\CA5\part 2\one\DFlipFlop / module Pad_Bond / page Page0 
.ENDS

.SUBCKT PadBidirHE_2.0u DataIn DataInB DataInUnBuf DataOut OE Pad Gnd Subs Vdd
MN_4_1 OEB OE Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MN_4_2 N29 DataOut Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MN_4_3 N20 OE N29 Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MN_4_4 N29 OEB Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MN_4_5 Pad N29 Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=10
MN_4_6 DataInB DataInUnBuf Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=2
MN_4_7 DataIn DataInB Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=4
XPad_Bond_1 Pad Subs Pad_Bond
* Page Size:  5x7
* S-Edit  Bidirectional Pad
* Designed by: D.Gunawan, J.Luo  Jan 12, 2025  14:21:54
* Schematic generated by S-Edit
* from file D:\Desktop\Electronic Digital\CA5\part 2\one\DFlipFlop / module PadBidirHE_2.0u / page Page0 
MP_4_1 OEB OE Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MP_4_2 N20 DataOut Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=2
MP_4_3 N29 OEB N20 Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=2
MP_4_4 N20 OE Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MP_4_5 Pad N20 Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=10
MP_4_6 DataInB DataInUnBuf Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=2
MP_4_7 DataIn DataInB Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=4
R1 Pad DataInUnBuf 100 TC1=0.0 TC2=0.0
.ENDS

.SUBCKT PadBidirHE DataIn DataInB DataInUnBuf DataOut OE Pad Gnd Subs Vdd
XPadBidirHE_2.0u_1 DataIn DataInB DataInUnBuf DataOut OE Pad Gnd Subs Vdd
+ PadBidirHE_2.0u
* Page Size:  5x7
* S-Edit  Bidirectional Pad
* Designed by: D.Gunawan, J.Luo  Jan 12, 2025  14:21:54
* Schematic generated by S-Edit
* from file D:\Desktop\Electronic Digital\CA5\part 2\one\DFlipFlop / module PadBidirHE / page Page0 
.ENDS

.SUBCKT PadInC DataIn DataInB DataInUnBuf Pad Gnd Subs Vdd
XPadBidirHE_1 DataIn DataInB DataInUnBuf Gnd Gnd Pad Gnd Subs Vdd PadBidirHE
* Page Size:  5x7
* S-Edit  Input Pad
* Designed by: D.Gunawan, J.Luo  Jan 12, 2025  14:20:40
* Schematic generated by S-Edit
* from file D:\Desktop\Electronic Digital\CA5\part 2\one\DFlipFlop / module PadInC / page Page0 
.ENDS

.SUBCKT NAND2 A B Out Gnd Vdd
M3 Out B 1 Gnd NMOS W='28*l' L='2*l' AS='148*l*l' AD='84*l*l' PS='68*l' PD='34*l' M=1
M4 1 A Gnd Gnd NMOS W='28*l' L='2*l' AS='84*l*l' AD='144*l*l' PS='34*l' PD='68*l' M=1
* Page Size:  5x7
* S-Edit  2-Input NAND Gate (TIB)
* Designed by: J. Luo  Jan 12, 2025  14:18:33
* Schematic generated by S-Edit
* from file D:\Desktop\Electronic Digital\CA5\part 2\one\DFlipFlop / module NAND2 / page Page0 
M2 Out B Vdd Vdd PMOS W='28*l' L='2*l' AS='144*l*l' AD='84*l*l' PS='68*l' PD='34*l' M=1
M1 Out A Vdd Vdd PMOS W='28*l' L='2*l' AS='84*l*l' AD='144*l*l' PS='34*l' PD='68*l' M=1
.ENDS

.SUBCKT NAND3 A B C Out Gnd Vdd
M4 Out C 1 Gnd NMOS W='28*l' L='2*l' AS='148*l*l' AD='84*l*l' PS='68*l' PD='34*l' M=1
M5 1 B 2 Gnd NMOS W='28*l' L='2*l' AS='84*l*l' AD='84*l*l' PS='34*l' PD='34*l' M=1
M6 2 A Gnd Gnd NMOS W='28*l' L='2*l' AS='84*l*l' AD='144*l*l' PS='34*l' PD='68*l' M=1
* Page Size:  5x7
* S-Edit  3-Input NAND Gate (TIB)
* Designed by: J. Luo   Jan 12, 2025  14:18:33
* Schematic generated by S-Edit
* from file D:\Desktop\Electronic Digital\CA5\part 2\one\DFlipFlop / module NAND3 / page Page0 
M1 Out A Vdd Vdd PMOS W='28*l' L='2*l' AS='84*l*l' AD='144*l*l' PS='34*l' PD='68*l' M=1
M2 Out B Vdd Vdd PMOS W='28*l' L='2*l' AS='84*l*l' AD='84*l*l' PS='34*l' PD='34*l' M=1
M3 Out C Vdd Vdd PMOS W='28*l' L='2*l' AS='148*l*l' AD='84*l*l' PS='68*l' PD='34*l' M=1
.ENDS

.SUBCKT D_flip_flop clk D Q Gnd Vdd
XNAND2_3 N7 N8 Q Gnd Vdd NAND2
XNAND2_4 Q N13 N8 Gnd Vdd NAND2
XNAND2_5 N11 N7 N17 Gnd Vdd NAND2
XNAND2_6 N17 clk N7 Gnd Vdd NAND2
XNAND2_7 N13 D N11 Gnd Vdd NAND2
XNAND3_1 N7 clk N11 N13 Gnd Vdd NAND3
.ENDS

.SUBCKT PadOut DataOut Pad Gnd Subs Vdd
XPadBidirHE_1 N6 N5 N4 DataOut Vdd Pad Gnd Subs Vdd PadBidirHE
* Page Size:  5x7
* S-Edit  Output Pad
* Designed by: D.Gunawan, J.Luo  Jan 12, 2025  14:21:54
* Schematic generated by S-Edit
* from file D:\Desktop\Electronic Digital\CA5\part 2\one\DFlipFlop / module PadOut / page Page0 
.ENDS

* Main circuit: shift_register_4bbit
XD_flip_flop_1 clk N4 N11 Gnd Vdd D_flip_flop
XD_flip_flop_2 clk N11 N9 Gnd Vdd D_flip_flop
XD_flip_flop_3 clk N9 N6 Gnd Vdd D_flip_flop
XD_flip_flop_4 clk N6 N5 Gnd Vdd D_flip_flop
XPadInC_1 N4 N3 N2 in Gnd Subs Vdd PadInC
XPadOut_1 N5 out Gnd Subs Vdd PadOut
* End of main circuit: shift_register_4bbit
